`define DATA_BITS 32
`define ADDR_BITS 32
`define BRANCH_CTRL_BITS 2
`define IMM_TYPE 3
`define REG_ADDR 5
`define OPCODE_BITS 7
`define BRANCH_TYPE_BITS 2
`define ALU_TYPE_BITS 3
`define FUNCT3_BITS 3
`define FUNCT7_BITS 7
`define FORWARDMUX 2
`define ALU_CTRL_BITS 5
`define INSTR_COUNT_TYPES 2
`define COUNTER_BITS 64
`define CSR_IMM_BITS 12
`define MUL_BITS 64

