`define CPU_CYCLE     11.5 // 100Mhz
`define MAX           9000000 // 3000000
`define AXI_CYCLE     25.0 // 40Mhz